version https://git-lfs.github.com/spec/v1
oid sha256:ec7a929d818dd4b8fdcb00054c67882e5c2217619e659e1ab82670338955f105
size 184
